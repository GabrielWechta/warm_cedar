LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE pack IS

	FUNCTION nextCRC
	(
		data : STD_LOGIC_VECTOR(7 DOWNTO 0);
		prevCRC : STD_LOGIC_VECTOR(7 DOWNTO 0)
	) RETURN STD_LOGIC_VECTOR;

END pack;

PACKAGE BODY pack IS

	FUNCTION nextCRC
	(
		data : STD_LOGIC_VECTOR(7 DOWNTO 0);
		prevCRC : STD_LOGIC_VECTOR(7 DOWNTO 0)
	)
		RETURN STD_LOGIC_VECTOR IS

		VARIABLE D : STD_LOGIC_VECTOR(7 DOWNTO 0);
		VARIABLE C : STD_LOGIC_VECTOR(7 DOWNTO 0);
		VARIABLE newCRC : STD_LOGIC_VECTOR(7 DOWNTO 0);

	BEGIN
		D := data;
		C := prevCRC;

		newCRC(0) := D(7) XOR D(6) XOR D(0) XOR C(0) XOR C(6) XOR C(7);
		newCRC(1) := D(6) XOR D(1) XOR D(0) XOR C(0) XOR C(1) XOR C(6);
		newCRC(2) := D(6) XOR D(2) XOR D(1) XOR D(0) XOR C(0) XOR C(1)
		XOR C(2) XOR C(6);
		newCRC(3) := D(7) XOR D(3) XOR D(2) XOR D(1) XOR C(1) XOR C(2)
		XOR C(3) XOR C(7);
		newCRC(4) := D(4) XOR D(3) XOR D(2) XOR C(2) XOR C(3) XOR C(4);
		newCRC(5) := D(5) XOR D(4) XOR D(3) XOR C(3) XOR C(4) XOR C(5);
		newCRC(6) := D(6) XOR D(5) XOR D(4) XOR C(4) XOR C(5) XOR C(6);
		newCRC(7) := D(7) XOR D(6) XOR D(5) XOR C(5) XOR C(6) XOR C(7);

		RETURN newCRC;
	END nextCRC;

END pack;